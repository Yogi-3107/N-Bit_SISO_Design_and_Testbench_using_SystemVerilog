interface intf #(parameter N = 4) (input logic clk);
  logic rst;
  logic serial_in;
  logic serial_out;
endinterface